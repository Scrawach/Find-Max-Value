// ----------
// TIME SCALE
// ----------

`timescale 1ns / 1ns
